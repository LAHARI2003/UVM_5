// This is DIMC TILE wrap env class instantiating feature_buffer_env, kernel_mem_env, 
// output_buffer_env, psin_env, addin_env, register_env (replaces computation_env), 
// p18_dimc_tile_wrap_virtual_sequencer

class p18_dimc_tile_wrap_env extends uvm_env;

  // Sub-environment instances
  istream_env#(64) m_feature_buffer_env;
  virtual istream_if#(64) vif;

  dpmem_env#(64,9)     m_kernel_mem_env;
  virtual dpmem_if#(64,9) kernel_mem_vif;

  ostream_env#(64)  m_output_buffer_env;
  virtual ostream_if#(64) ostream_vif;

  //psin_env           m_psin_env;
  istream_env#(32)   m_psin_env;
  virtual istream_if#(32) psin_vif;

  spmem_env#(64,4)          m_addin_env;
  virtual spmem_if#(64,4)   addin_vif;

  // New register_env replaces computation_env
  register_env    m_register_env;
  virtual register_if register_vif;

  p18_dimc_tile_wrap_virtual_sequencer  v_seqr;

  p18_dimc_tile_wrap_scoreboard#(64) dimc_tile_wrap_scoreboard;

  `uvm_component_utils(p18_dimc_tile_wrap_env)

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    // Create sub-environments
    m_feature_buffer_env = istream_env#(64)::type_id::create("m_feature_buffer_env", this);
    m_kernel_mem_env     = dpmem_env#(64,9)::type_id::create("m_kernel_mem_env", this);
    m_output_buffer_env  = ostream_env#(64)::type_id::create("m_output_buffer_env", this);
    m_psin_env           = istream_env#(32)::type_id::create("m_psin_env", this);
    m_addin_env          = spmem_env#(64,4)::type_id::create("m_addin_env", this);
    // Create register_env instead of computation_env
    m_register_env       = register_env::type_id::create("m_register_env", this);
    
 
    v_seqr               = p18_dimc_tile_wrap_virtual_sequencer::type_id::create("v_seqr", this);
    dimc_tile_wrap_scoreboard = p18_dimc_tile_wrap_scoreboard#(64)::type_id::create("dimc_tile_wrap_scoreboard", this);

   if (!uvm_config_db#(virtual istream_if#(64))::get(this, "*", "feature_buffer_vif", vif))
      `uvm_fatal("NOVIF", "Virtual interface must be set for vif")

   if (!uvm_config_db#(virtual istream_if#(32))::get(this, "*", "psin_vif", psin_vif))
      `uvm_fatal("NOVIF", "Virtual interface must be set for psin_vif")

   if (!uvm_config_db#(virtual ostream_if#(64))::get(this, "", "ostream_vif", ostream_vif))
      `uvm_fatal("NOVIF", "Virtual interface must be set for ostream_vif")

   if (!uvm_config_db#(virtual spmem_if#(64,4))::get(this, "", "addin_vif", addin_vif))
      `uvm_fatal("NOVIF", "Virtual interface must be set for addin_vif")

  if (!uvm_config_db#(virtual dpmem_if#(64,9))::get(this, "", "kernel_mem_vif", kernel_mem_vif))
      `uvm_fatal("NOVIF", "Virtual interface must be set for kernel_mem_vif") 

  // Get register_vif instead of computation_vif
  if (!uvm_config_db#(virtual register_if)::get(this, "", "register_vif", register_vif))
      `uvm_fatal("NOVIF", "Virtual interface must be set for register_vif")

endfunction

  // Add connect_phase or other phases as needed
       function void connect_phase(uvm_phase phase);
    		super.connect_phase(phase);
    		v_seqr.seqr_feature_buffer		= m_feature_buffer_env.m_agent.m_sequencer;		//sequencer kmem axi
    		v_seqr.seqr_kernel_mem  		= m_kernel_mem_env.m_agent.m_sequencer;	 	
    		v_seqr.seqr_output_buffer        	= m_output_buffer_env.m_agent.m_sequencer;		

		v_seqr.seqr_psin			= m_psin_env.m_agent.m_sequencer;		
		v_seqr.seqr_addin			= m_addin_env.m_agent.m_sequencer;
                // Connect register sequencer instead of computation sequencer
                v_seqr.seqr_register                    = m_register_env.m_agent.m_sequencer;

                m_feature_buffer_env.m_agent.vif                 = vif;
                m_feature_buffer_env.m_agent.m_driver.vif        = vif;
                m_feature_buffer_env.m_agent.m_monitor.vif        = vif;

                m_psin_env.m_agent.vif                  = psin_vif;
                m_psin_env.m_agent.m_driver.vif         = psin_vif;
                m_psin_env.m_agent.m_monitor.vif        = psin_vif;

                m_addin_env.m_agent.vif                 = addin_vif;
                m_addin_env.m_agent.m_driver.vif        = addin_vif;

                m_output_buffer_env.m_agent.m_driver.vif = ostream_vif;
               	m_output_buffer_env.m_agent.m_sequencer.vif = ostream_vif;
                m_output_buffer_env.m_agent.m_monitor.vif = ostream_vif;
                m_output_buffer_env.m_agent.m_monitor.ostream_rd_port.connect(dimc_tile_wrap_scoreboard.imp_ostream_rd_port);

                m_kernel_mem_env.m_agent.vif                 = kernel_mem_vif;
                m_kernel_mem_env.m_agent.m_driver.vif        = kernel_mem_vif;

                // Connect register interface to register agent and driver
                m_register_env.m_agent.vif                   = register_vif;
                m_register_env.m_agent.m_driver.vif          = register_vif;

  	endfunction


endclass
