// This istream_directed_write_sequence generated istream_seq_item 16 times
// and pass it to the istream_sequencer 
// This reads the input frame from the file istream_data_unique_64x16.txt and
// saves it into the istream_data_ip of two dimensional array of 16 rows and 64
// columns
// This stores istream_data_ip row gets driven to req.istream_data field
class istream_directed_random_burst_write_sequence #(int DATA_WIDTH = 32) extends uvm_sequence #(istream_seq_item);

  `uvm_object_utils(istream_directed_random_burst_write_sequence#(DATA_WIDTH))
  //`uvm_param_utils(feature_directed_write_sequence#(DATA_WIDTH))

  function new(string name = "istream_directed_random_burst_write_sequence");
    super.new(name);
  endfunction

  logic [DATA_WIDTH-1:0] istream_data_ip [];
  int i;
  int size;
  int k=0;
  int l=0;
  int j =0;
  string file_path;

 
  istream_seq_item#(DATA_WIDTH) req;
  ip_stall_rand	 tr_stall_rand;

  task body();
   begin
    istream_data_ip = new[size];
    //$readmemh("./input_data/feature_data_unique_64x16.txt", feat_data_ip) ;
    $readmemh(file_path, istream_data_ip) ;
    

    for(i = 0; i<size; i++)
      begin : istream_wr

        tr_stall_rand	= ip_stall_rand::type_id::create("tr_stall_rand");
        //assert(req.randomize());
	tr_stall_rand.randomize();
        $display("burst_len = %0d; inter_burst_latency = %0d \n time = %0g", tr_stall_rand.burst_len,tr_stall_rand.inter_bus_latency,$time);

       if ( tr_stall_rand.burst_len > (size-i) ) begin
         tr_stall_rand.burst_len = size-i;
       end
       for(k = 0; k<tr_stall_rand.burst_len; k++)
	   begin
		req = istream_seq_item#(DATA_WIDTH)::type_id::create("req");
                req.istream_valid = 1'b1;
                req.istream_data  = istream_data_ip[j];
		j=j+1;
                // `uvm_do_with(req,{req.feat_valid==1'b1;req.feat_data  == feat_data_ip[i];});
                start_item(req);
                finish_item(req);
          end
        
       for(l = 0; l<tr_stall_rand.inter_bus_latency; l++)
	  begin
	        req = istream_seq_item#(DATA_WIDTH)::type_id::create("req");
                req.istream_valid = 1'b0;
                req.istream_data  = 0;
	        // `uvm_do_with(req,{req.feat_valid==1'b1;req.feat_data  == feat_data_ip[i];});
                start_item(req);
                finish_item(req);
         end

        i = i+tr_stall_rand.burst_len-1;   
 
     end : istream_wr

 // Disabling istream buffer
        req.istream_valid = 1'b0;
        req.istream_data  = 64'h0;

        //`uvm_do_with(req,{req.feat_valid==1'b0;req.feat_data  == 64'h0;});

       //`uvm_do(req);
        start_item(req);
        finish_item(req);

    end
  endtask

endclass
